/*
	this is my first and gate.
*/
module And_Gate(A, B, F);

	input A, B;
	output F;
		wire A, B;
		wire F;
		
		assign F = A & B;

endmodule